architecture arch of seven_segment_control is
signal r_reg, r_next : unsigned (COUNTER_BITS-1 downto 0) := (others=> '0');
signal num : STD_LOGIC_VECTOR(3 downto 0);
signal counter : STD_LOGIC_VECTOR(COUNTER_BITS-1 downto 0);
signal an_sel : STD_LOGIC_VECTOR(1 downto 0);

begin
an_sel <= counter(COUNTER_BITS-1 downto COUNTER_BITS-2);
--selected signal assignment statement for seven segment display
with num select
seg(6 downto 0) <= "1000000" when "0000",--0
"1111001" when "0001",--1
"0100100" when "0010",--2
"0110000" when "0011",--3
"0011001" when "0100",--4
"0010010" when "0101",--5
"0000010" when "0110",--6
"1111000" when "0111",--7
"0000000" when "1000",--8
"0010000" when "1001",--9
"0001000" when "1010",--A
"0000011" when "1011",--B
"1000110" when "1100",--C
"0100001" when "1101",--D
"0000110" when "1110",--E
"0001110" when others;--F



--mux with input btn(1 downto 0) 
with an_sel select
num <= data_in(3 downto 0) when "00",
data_in(7 downto 4) when "01",
data_in(11 downto 8) when "10",
data_in(15 downto 12) when others;

--decimal point logic
with an_sel select
dp <= not dp_in(0) when "00",
not dp_in(1) when "01",
not dp_in(2) when "10",
not dp_in(3) when others;

--anode logic 
an <= "111" & blank(0) when (an_sel = "00") else
"11" & blank(1) & '1' when (an_sel = "01") else
'1' & blank(2) & "11" when (an_sel = "10") else
blank(3) & "111";


process(clk)
begin
if clk'event and clk = '1' then
r_reg <= r_next;
end if;

end process;
r_next <= r_reg+1;
counter <= std_logic_vector(r_reg);
end arch;